module mesh_twoxone(rt_clk, neu_clk, rt_reset, neu_reset,
                    north_out_1_1, north_out_1_2, south_out_1_1, south_out_1_2,
                    west_out_1_1,
                    north_in_1_1, north_in_1_2, south_in_1_1, south_in_1_2,
                    west_in_1_1,
                    write_en_north_1_1, write_en_north_1_2, write_en_south_1_1, write_en_south_1_2,
                    write_en_west_1_1,
                    write_req_);

